module AC(
	


);
